ENTITY mux_2x1_Wbits IS
GENERIC (W : NATURAL := 16);
